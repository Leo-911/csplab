`ifndef DATA_TYPE_SVH_
`define DATA_TYPE_SVH_
// I/O types
typedef logic signed [15:0] r_t;
typedef logic signed [7:0]  rho_t;
typedef logic signed [20:0] eps_t;
typedef logic [7:0]         theta_t;

// Port types
typedef logic signed [15:0] phi_t;
typedef logic signed [15:0] gamma_t;
typedef logic signed [15:0] mag_t;
typedef logic signed [12:0] ang_t;
typedef logic signed [15:0] lambda_t;

// Internal types
typedef logic signed [11:0] ambm_t;
typedef logic [9:0]         PI_t;
typedef logic [7:0]         ratio_t;

`endif // DATA_TYPE_SVH_
